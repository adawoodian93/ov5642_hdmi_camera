`timescale 1ns / 1ps
module ov5642_init_regs (
  input wire [9:0]  i_addr,
  output reg [23:0] o_data, //[23:8] = addr; [7:0] = data
  output reg        o_verify
);

  always @(*) begin
    case (i_addr)
      10'd0: {o_verify, o_data} <= {1'b1, 24'h3103_93};
      10'd1: {o_verify, o_data} <= {1'b1, 24'h3008_82};
      /*10'd2: {o_verify, o_data} <= {1'b1, 24'h3017_7f};
      10'd3: {o_verify, o_data} <= {1'b1, 24'h3018_fc};
      10'd4: {o_verify, o_data} <= {1'b1, 24'h3810_c2};
      10'd5: {o_verify, o_data} <= {1'b1, 24'h3615_f0};
      10'd6: {o_verify, o_data} <= {1'b1, 24'h3000_00};
      10'd7: {o_verify, o_data} <= {1'b1, 24'h3001_00};
      10'd8: {o_verify, o_data} <= {1'b1, 24'h3002_00};
      10'd9: {o_verify, o_data} <= {1'b1, 24'h3003_00};
      10'd10: {o_verify, o_data} <= {1'b1, 24'h3004_ff};
      10'd11: {o_verify, o_data} <= {1'b1, 24'h3030_2b};
      10'd12: {o_verify, o_data} <= {1'b1, 24'h3011_08};
      10'd13: {o_verify, o_data} <= {1'b1, 24'h3010_10};
      10'd14: {o_verify, o_data} <= {1'b1, 24'h3604_60};
      10'd15: {o_verify, o_data} <= {1'b1, 24'h3622_60};
      10'd16: {o_verify, o_data} <= {1'b1, 24'h3621_09};
      10'd17: {o_verify, o_data} <= {1'b1, 24'h3709_00};
      10'd18: {o_verify, o_data} <= {1'b1, 24'h4000_21};
      10'd19: {o_verify, o_data} <= {1'b1, 24'h401d_22};
      10'd20: {o_verify, o_data} <= {1'b1, 24'h3600_54};
      10'd21: {o_verify, o_data} <= {1'b1, 24'h3605_04};
      10'd22: {o_verify, o_data} <= {1'b1, 24'h3606_3f};
      10'd23: {o_verify, o_data} <= {1'b1, 24'h3c01_80};
      10'd24: {o_verify, o_data} <= {1'b1, 24'h300d_22};
      10'd25: {o_verify, o_data} <= {1'b1, 24'h3623_22};
      10'd26: {o_verify, o_data} <= {1'b1, 24'h5000_4f};
      10'd27: {o_verify, o_data} <= {1'b1, 24'h5020_04};
      10'd28: {o_verify, o_data} <= {1'b1, 24'h5181_79};
      10'd29: {o_verify, o_data} <= {1'b1, 24'h5182_00};
      10'd30: {o_verify, o_data} <= {1'b1, 24'h5185_22};
      10'd31: {o_verify, o_data} <= {1'b1, 24'h5197_01};
      10'd32: {o_verify, o_data} <= {1'b1, 24'h5500_0a};
      10'd33: {o_verify, o_data} <= {1'b1, 24'h5504_00};
      10'd34: {o_verify, o_data} <= {1'b1, 24'h5505_7f};
      10'd35: {o_verify, o_data} <= {1'b1, 24'h5080_08};
      10'd36: {o_verify, o_data} <= {1'b1, 24'h300e_18};
      10'd37: {o_verify, o_data} <= {1'b1, 24'h4610_00};
      10'd38: {o_verify, o_data} <= {1'b1, 24'h471d_05};
      10'd39: {o_verify, o_data} <= {1'b1, 24'h4708_06};
      10'd40: {o_verify, o_data} <= {1'b1, 24'h370c_a0};
      10'd41: {o_verify, o_data} <= {1'b1, 24'h3808_0a};
      10'd42: {o_verify, o_data} <= {1'b1, 24'h3809_20};
      10'd43: {o_verify, o_data} <= {1'b1, 24'h380a_07};
      10'd44: {o_verify, o_data} <= {1'b1, 24'h380b_98};
      10'd45: {o_verify, o_data} <= {1'b1, 24'h380c_0c};
      10'd46: {o_verify, o_data} <= {1'b1, 24'h380d_80};
      10'd47: {o_verify, o_data} <= {1'b1, 24'h380e_07};
      10'd48: {o_verify, o_data} <= {1'b1, 24'h380f_d0};
      10'd49: {o_verify, o_data} <= {1'b1, 24'h5687_94};
      10'd50: {o_verify, o_data} <= {1'b1, 24'h501f_00};
      10'd51: {o_verify, o_data} <= {1'b1, 24'h5000_4f};
      10'd52: {o_verify, o_data} <= {1'b1, 24'h5001_cf};
      10'd53: {o_verify, o_data} <= {1'b1, 24'h4300_61}; //format control register RGB565
      10'd54: {o_verify, o_data} <= {1'b1, 24'h4300_61}; //format control register RGB565
      10'd55: {o_verify, o_data} <= {1'b1, 24'h460b_35};
      10'd56: {o_verify, o_data} <= {1'b1, 24'h471d_00};
      10'd57: {o_verify, o_data} <= {1'b1, 24'h3002_0c};
      10'd58: {o_verify, o_data} <= {1'b1, 24'h3002_00};
      10'd59: {o_verify, o_data} <= {1'b1, 24'h4713_03};
      10'd60: {o_verify, o_data} <= {1'b1, 24'h471c_50};
      10'd61: {o_verify, o_data} <= {1'b1, 24'h4721_02};
      10'd62: {o_verify, o_data} <= {1'b1, 24'h4402_90};
      10'd63: {o_verify, o_data} <= {1'b1, 24'h460c_22};
      10'd64: {o_verify, o_data} <= {1'b1, 24'h3815_44};
      10'd65: {o_verify, o_data} <= {1'b1, 24'h3503_07};
      10'd66: {o_verify, o_data} <= {1'b1, 24'h3501_73};
      10'd67: {o_verify, o_data} <= {1'b1, 24'h3502_80};
      10'd68: {o_verify, o_data} <= {1'b1, 24'h350b_00};
      10'd69: {o_verify, o_data} <= {1'b1, 24'h3818_c8};
      10'd70: {o_verify, o_data} <= {1'b1, 24'h3801_88};
      10'd71: {o_verify, o_data} <= {1'b1, 24'h3824_11};
      10'd72: {o_verify, o_data} <= {1'b1, 24'h3a00_78};
      10'd73: {o_verify, o_data} <= {1'b1, 24'h3a1a_04};
      10'd74: {o_verify, o_data} <= {1'b1, 24'h3a13_30};
      10'd75: {o_verify, o_data} <= {1'b1, 24'h3a18_00};
      10'd76: {o_verify, o_data} <= {1'b1, 24'h3a19_7c};
      10'd77: {o_verify, o_data} <= {1'b1, 24'h3a08_12};
      10'd78: {o_verify, o_data} <= {1'b1, 24'h3a09_c0};
      10'd79: {o_verify, o_data} <= {1'b1, 24'h3a0a_0f};
      10'd80: {o_verify, o_data} <= {1'b1, 24'h3a0b_a0};
      10'd81: {o_verify, o_data} <= {1'b1, 24'h350c_07};
      10'd82: {o_verify, o_data} <= {1'b1, 24'h350d_d0};
      10'd83: {o_verify, o_data} <= {1'b1, 24'h3a0d_08};
      10'd84: {o_verify, o_data} <= {1'b1, 24'h3a0e_06};
      10'd85: {o_verify, o_data} <= {1'b1, 24'h3500_00};
      10'd86: {o_verify, o_data} <= {1'b1, 24'h3501_00};
      10'd87: {o_verify, o_data} <= {1'b1, 24'h3502_00};
      10'd88: {o_verify, o_data} <= {1'b1, 24'h350a_00};
      10'd89: {o_verify, o_data} <= {1'b1, 24'h350b_00};
      10'd90: {o_verify, o_data} <= {1'b1, 24'h3503_00};
      10'd91: {o_verify, o_data} <= {1'b1, 24'h3030_2b};
      10'd92: {o_verify, o_data} <= {1'b1, 24'h3a02_00};
      10'd93: {o_verify, o_data} <= {1'b1, 24'h3a03_7d};
      10'd94: {o_verify, o_data} <= {1'b1, 24'h3a04_00};
      10'd95: {o_verify, o_data} <= {1'b1, 24'h3a14_00};
      10'd96: {o_verify, o_data} <= {1'b1, 24'h3a15_7d};
      10'd97: {o_verify, o_data} <= {1'b1, 24'h3a16_00};
      10'd98: {o_verify, o_data} <= {1'b1, 24'h3a00_78};
      10'd99: {o_verify, o_data} <= {1'b1, 24'h3a08_09};
      10'd100: {o_verify, o_data} <= {1'b1, 24'h3a09_60};
      10'd101: {o_verify, o_data} <= {1'b1, 24'h3a0a_07};
      10'd102: {o_verify, o_data} <= {1'b1, 24'h3a0b_d0};
      10'd103: {o_verify, o_data} <= {1'b1, 24'h3a0d_10};
      10'd104: {o_verify, o_data} <= {1'b1, 24'h3a0e_0d};
      10'd105: {o_verify, o_data} <= {1'b1, 24'h4407_04};
      10'd106: {o_verify, o_data} <= {1'b1, 24'h5193_70};
      10'd107: {o_verify, o_data} <= {1'b1, 24'h589b_00};
      10'd108: {o_verify, o_data} <= {1'b1, 24'h589a_c0};
      10'd109: {o_verify, o_data} <= {1'b1, 24'h401e_20};
      10'd110: {o_verify, o_data} <= {1'b1, 24'h4001_42};
      10'd111: {o_verify, o_data} <= {1'b1, 24'h401c_06};
      10'd112: {o_verify, o_data} <= {1'b1, 24'h3825_ac};
      10'd113: {o_verify, o_data} <= {1'b1, 24'h3827_0c};
      10'd114: {o_verify, o_data} <= {1'b1, 24'h5402_3f};
      10'd115: {o_verify, o_data} <= {1'b1, 24'h5403_00};
      10'd116: {o_verify, o_data} <= {1'b1, 24'h3406_00};
      10'd117: {o_verify, o_data} <= {1'b1, 24'h5180_ff};
      10'd118: {o_verify, o_data} <= {1'b1, 24'h5181_52};
      10'd119: {o_verify, o_data} <= {1'b1, 24'h5182_11};
      10'd120: {o_verify, o_data} <= {1'b1, 24'h5183_14};
      10'd121: {o_verify, o_data} <= {1'b1, 24'h5184_25};
      10'd122: {o_verify, o_data} <= {1'b1, 24'h5185_24};
      10'd123: {o_verify, o_data} <= {1'b1, 24'h5186_06};
      10'd124: {o_verify, o_data} <= {1'b1, 24'h5187_08};
      10'd125: {o_verify, o_data} <= {1'b1, 24'h5188_08};
      10'd126: {o_verify, o_data} <= {1'b1, 24'h5189_7c};
      10'd127: {o_verify, o_data} <= {1'b1, 24'h518a_60};
      10'd128: {o_verify, o_data} <= {1'b1, 24'h518b_b2};
      10'd129: {o_verify, o_data} <= {1'b1, 24'h518c_b2};
      10'd130: {o_verify, o_data} <= {1'b1, 24'h518d_44};
      10'd131: {o_verify, o_data} <= {1'b1, 24'h518e_3d};
      10'd132: {o_verify, o_data} <= {1'b1, 24'h518f_58};
      10'd133: {o_verify, o_data} <= {1'b1, 24'h5190_46};
      10'd134: {o_verify, o_data} <= {1'b1, 24'h5191_f8};
      10'd135: {o_verify, o_data} <= {1'b1, 24'h5192_04};
      10'd136: {o_verify, o_data} <= {1'b1, 24'h5193_70};
      10'd137: {o_verify, o_data} <= {1'b1, 24'h5194_f0};
      10'd138: {o_verify, o_data} <= {1'b1, 24'h5195_f0};
      10'd139: {o_verify, o_data} <= {1'b1, 24'h5196_03};
      10'd140: {o_verify, o_data} <= {1'b1, 24'h5197_01};
      10'd141: {o_verify, o_data} <= {1'b1, 24'h5198_04};
      10'd142: {o_verify, o_data} <= {1'b1, 24'h5199_12};
      10'd143: {o_verify, o_data} <= {1'b1, 24'h519a_04};
      10'd144: {o_verify, o_data} <= {1'b1, 24'h519b_00};
      10'd145: {o_verify, o_data} <= {1'b1, 24'h519c_06};
      10'd146: {o_verify, o_data} <= {1'b1, 24'h519d_82};
      10'd147: {o_verify, o_data} <= {1'b1, 24'h519e_00};
      10'd148: {o_verify, o_data} <= {1'b1, 24'h5025_80};
      10'd149: {o_verify, o_data} <= {1'b1, 24'h5583_40};
      10'd150: {o_verify, o_data} <= {1'b1, 24'h5584_40};
      10'd151: {o_verify, o_data} <= {1'b1, 24'h5580_02};
      10'd152: {o_verify, o_data} <= {1'b1, 24'h5000_cf};
      10'd153: {o_verify, o_data} <= {1'b1, 24'h3710_10};
      10'd154: {o_verify, o_data} <= {1'b1, 24'h3632_51};
      10'd155: {o_verify, o_data} <= {1'b1, 24'h3702_10};
      10'd156: {o_verify, o_data} <= {1'b1, 24'h3703_b2};
      10'd157: {o_verify, o_data} <= {1'b1, 24'h3704_18};
      10'd158: {o_verify, o_data} <= {1'b1, 24'h370b_40};
      10'd159: {o_verify, o_data} <= {1'b1, 24'h370d_03};
      10'd160: {o_verify, o_data} <= {1'b1, 24'h3631_01};
      10'd161: {o_verify, o_data} <= {1'b1, 24'h3632_52};
      10'd162: {o_verify, o_data} <= {1'b1, 24'h3606_24};
      10'd163: {o_verify, o_data} <= {1'b1, 24'h3620_96};
      10'd164: {o_verify, o_data} <= {1'b1, 24'h5785_07};
      10'd165: {o_verify, o_data} <= {1'b1, 24'h3a13_30};
      10'd166: {o_verify, o_data} <= {1'b1, 24'h3600_52};
      10'd167: {o_verify, o_data} <= {1'b1, 24'h3604_48};
      10'd168: {o_verify, o_data} <= {1'b1, 24'h3606_1b};
      10'd169: {o_verify, o_data} <= {1'b1, 24'h370d_0b};
      10'd170: {o_verify, o_data} <= {1'b1, 24'h370f_c0};
      10'd171: {o_verify, o_data} <= {1'b1, 24'h3709_01};
      10'd172: {o_verify, o_data} <= {1'b1, 24'h3823_00};
      10'd173: {o_verify, o_data} <= {1'b1, 24'h5007_00};
      10'd174: {o_verify, o_data} <= {1'b1, 24'h5009_00};
      10'd175: {o_verify, o_data} <= {1'b1, 24'h5011_00};
      10'd176: {o_verify, o_data} <= {1'b1, 24'h5013_00};
      10'd177: {o_verify, o_data} <= {1'b1, 24'h519e_00};
      10'd178: {o_verify, o_data} <= {1'b1, 24'h5086_00};
      10'd179: {o_verify, o_data} <= {1'b1, 24'h5087_00};
      10'd180: {o_verify, o_data} <= {1'b1, 24'h5088_00};
      10'd181: {o_verify, o_data} <= {1'b1, 24'h5089_00};
      10'd182: {o_verify, o_data} <= {1'b1, 24'h302b_00};
      10'd183: {o_verify, o_data} <= {1'b1, 24'h3503_07};
      10'd184: {o_verify, o_data} <= {1'b1, 24'h3011_07};
      10'd185: {o_verify, o_data} <= {1'b1, 24'h350c_04};
      10'd186: {o_verify, o_data} <= {1'b1, 24'h350d_58};
      10'd187: {o_verify, o_data} <= {1'b1, 24'h3801_8a};
      10'd188: {o_verify, o_data} <= {1'b1, 24'h3803_0a};
      10'd189: {o_verify, o_data} <= {1'b1, 24'h3804_07};
      10'd190: {o_verify, o_data} <= {1'b1, 24'h3805_80};
      10'd191: {o_verify, o_data} <= {1'b1, 24'h3806_04};
      10'd192: {o_verify, o_data} <= {1'b1, 24'h3807_38};
      10'd193: {o_verify, o_data} <= {1'b1, 24'h3808_07};
      10'd194: {o_verify, o_data} <= {1'b1, 24'h3809_80};
      10'd195: {o_verify, o_data} <= {1'b1, 24'h380a_04};
      10'd196: {o_verify, o_data} <= {1'b1, 24'h380b_38};
      10'd197: {o_verify, o_data} <= {1'b1, 24'h380c_09};
      10'd198: {o_verify, o_data} <= {1'b1, 24'h380d_d6};
      10'd199: {o_verify, o_data} <= {1'b1, 24'h380e_04};
      10'd200: {o_verify, o_data} <= {1'b1, 24'h380f_58};
      10'd201: {o_verify, o_data} <= {1'b1, 24'h381c_11};
      10'd202: {o_verify, o_data} <= {1'b1, 24'h381d_ba};
      10'd203: {o_verify, o_data} <= {1'b1, 24'h381e_04};
      10'd204: {o_verify, o_data} <= {1'b1, 24'h381f_48};
      10'd205: {o_verify, o_data} <= {1'b1, 24'h3820_04};
      10'd206: {o_verify, o_data} <= {1'b1, 24'h3821_18};
      10'd207: {o_verify, o_data} <= {1'b1, 24'h3a08_14};
      10'd208: {o_verify, o_data} <= {1'b1, 24'h3a09_e0};
      10'd209: {o_verify, o_data} <= {1'b1, 24'h3a0a_11};
      10'd210: {o_verify, o_data} <= {1'b1, 24'h3a0b_60};
      10'd211: {o_verify, o_data} <= {1'b1, 24'h3a0d_04};
      10'd212: {o_verify, o_data} <= {1'b1, 24'h3a0e_03};
      10'd213: {o_verify, o_data} <= {1'b1, 24'h5682_07};
      10'd214: {o_verify, o_data} <= {1'b1, 24'h5683_60};
      10'd215: {o_verify, o_data} <= {1'b1, 24'h5686_04};
      10'd216: {o_verify, o_data} <= {1'b1, 24'h5687_1c};
      10'd217: {o_verify, o_data} <= {1'b1, 24'h5001_7f};
      10'd218: {o_verify, o_data} <= {1'b1, 24'h3503_00};
      10'd219: {o_verify, o_data} <= {1'b1, 24'h3010_10};
      10'd220: {o_verify, o_data} <= {1'b1, 24'h5001_ff};
      10'd221: {o_verify, o_data} <= {1'b1, 24'h5583_50};
      10'd222: {o_verify, o_data} <= {1'b1, 24'h5584_50};
      10'd223: {o_verify, o_data} <= {1'b1, 24'h5580_02};
      10'd224: {o_verify, o_data} <= {1'b1, 24'h3c01_80};
      10'd225: {o_verify, o_data} <= {1'b1, 24'h3c00_04};
      10'd226: {o_verify, o_data} <= {1'b1, 24'h5800_48};
      10'd227: {o_verify, o_data} <= {1'b1, 24'h5801_31};
      10'd228: {o_verify, o_data} <= {1'b1, 24'h5802_21};
      10'd229: {o_verify, o_data} <= {1'b1, 24'h5803_1b};
      10'd230: {o_verify, o_data} <= {1'b1, 24'h5804_1a};
      10'd231: {o_verify, o_data} <= {1'b1, 24'h5805_1e};
      10'd232: {o_verify, o_data} <= {1'b1, 24'h5806_29};
      10'd233: {o_verify, o_data} <= {1'b1, 24'h5807_38};
      10'd234: {o_verify, o_data} <= {1'b1, 24'h5808_26};
      10'd235: {o_verify, o_data} <= {1'b1, 24'h5809_17};
      10'd236: {o_verify, o_data} <= {1'b1, 24'h580a_11};
      10'd237: {o_verify, o_data} <= {1'b1, 24'h580b_0e};
      10'd238: {o_verify, o_data} <= {1'b1, 24'h580c_0d};
      10'd239: {o_verify, o_data} <= {1'b1, 24'h580d_0e};
      10'd240: {o_verify, o_data} <= {1'b1, 24'h580e_13};
      10'd241: {o_verify, o_data} <= {1'b1, 24'h580f_1a};
      10'd242: {o_verify, o_data} <= {1'b1, 24'h5810_15};
      10'd243: {o_verify, o_data} <= {1'b1, 24'h5811_0d};
      10'd244: {o_verify, o_data} <= {1'b1, 24'h5812_08};
      10'd245: {o_verify, o_data} <= {1'b1, 24'h5813_05};
      10'd246: {o_verify, o_data} <= {1'b1, 24'h5814_04};
      10'd247: {o_verify, o_data} <= {1'b1, 24'h5815_05};
      10'd248: {o_verify, o_data} <= {1'b1, 24'h5816_09};
      10'd249: {o_verify, o_data} <= {1'b1, 24'h5817_0d};
      10'd250: {o_verify, o_data} <= {1'b1, 24'h5818_11};
      10'd251: {o_verify, o_data} <= {1'b1, 24'h5819_0a};
      10'd252: {o_verify, o_data} <= {1'b1, 24'h581a_04};
      10'd253: {o_verify, o_data} <= {1'b1, 24'h581b_00};
      10'd254: {o_verify, o_data} <= {1'b1, 24'h581c_00};
      10'd255: {o_verify, o_data} <= {1'b1, 24'h581d_01};
      10'd256: {o_verify, o_data} <= {1'b1, 24'h581e_06};
      10'd257: {o_verify, o_data} <= {1'b1, 24'h581f_09};
      10'd258: {o_verify, o_data} <= {1'b1, 24'h5820_12};
      10'd259: {o_verify, o_data} <= {1'b1, 24'h5821_0b};
      10'd260: {o_verify, o_data} <= {1'b1, 24'h5822_04};
      10'd261: {o_verify, o_data} <= {1'b1, 24'h5823_00};
      10'd262: {o_verify, o_data} <= {1'b1, 24'h5824_00};
      10'd263: {o_verify, o_data} <= {1'b1, 24'h5825_01};
      10'd264: {o_verify, o_data} <= {1'b1, 24'h5826_06};
      10'd265: {o_verify, o_data} <= {1'b1, 24'h5827_0a};
      10'd266: {o_verify, o_data} <= {1'b1, 24'h5828_17};
      10'd267: {o_verify, o_data} <= {1'b1, 24'h5829_0f};
      10'd268: {o_verify, o_data} <= {1'b1, 24'h582a_09};
      10'd269: {o_verify, o_data} <= {1'b1, 24'h582b_06};
      10'd270: {o_verify, o_data} <= {1'b1, 24'h582c_05};
      10'd271: {o_verify, o_data} <= {1'b1, 24'h582d_06};
      10'd272: {o_verify, o_data} <= {1'b1, 24'h582e_0a};
      10'd273: {o_verify, o_data} <= {1'b1, 24'h582f_0e};
      10'd274: {o_verify, o_data} <= {1'b1, 24'h5830_28};
      10'd275: {o_verify, o_data} <= {1'b1, 24'h5831_1a};
      10'd276: {o_verify, o_data} <= {1'b1, 24'h5832_11};
      10'd277: {o_verify, o_data} <= {1'b1, 24'h5833_0e};
      10'd278: {o_verify, o_data} <= {1'b1, 24'h5834_0e};
      10'd279: {o_verify, o_data} <= {1'b1, 24'h5835_0f};
      10'd280: {o_verify, o_data} <= {1'b1, 24'h5836_15};
      10'd281: {o_verify, o_data} <= {1'b1, 24'h5837_1d};
      10'd282: {o_verify, o_data} <= {1'b1, 24'h5838_6e};
      10'd283: {o_verify, o_data} <= {1'b1, 24'h5839_39};
      10'd284: {o_verify, o_data} <= {1'b1, 24'h583a_27};
      10'd285: {o_verify, o_data} <= {1'b1, 24'h583b_1f};
      10'd286: {o_verify, o_data} <= {1'b1, 24'h583c_1e};
      10'd287: {o_verify, o_data} <= {1'b1, 24'h583d_23};
      10'd288: {o_verify, o_data} <= {1'b1, 24'h583e_2f};
      10'd289: {o_verify, o_data} <= {1'b1, 24'h583f_41};
      10'd290: {o_verify, o_data} <= {1'b1, 24'h5840_0e};
      10'd291: {o_verify, o_data} <= {1'b1, 24'h5841_0c};
      10'd292: {o_verify, o_data} <= {1'b1, 24'h5842_0d};
      10'd293: {o_verify, o_data} <= {1'b1, 24'h5843_0c};
      10'd294: {o_verify, o_data} <= {1'b1, 24'h5844_0c};
      10'd295: {o_verify, o_data} <= {1'b1, 24'h5845_0c};
      10'd296: {o_verify, o_data} <= {1'b1, 24'h5846_0c};
      10'd297: {o_verify, o_data} <= {1'b1, 24'h5847_0c};
      10'd298: {o_verify, o_data} <= {1'b1, 24'h5848_0d};
      10'd299: {o_verify, o_data} <= {1'b1, 24'h5849_0e};
      10'd300: {o_verify, o_data} <= {1'b1, 24'h584a_0e};
      10'd301: {o_verify, o_data} <= {1'b1, 24'h584b_0a};
      10'd302: {o_verify, o_data} <= {1'b1, 24'h584c_0e};
      10'd303: {o_verify, o_data} <= {1'b1, 24'h584d_0e};
      10'd304: {o_verify, o_data} <= {1'b1, 24'h584e_10};
      10'd305: {o_verify, o_data} <= {1'b1, 24'h584f_10};
      10'd306: {o_verify, o_data} <= {1'b1, 24'h5850_11};
      10'd307: {o_verify, o_data} <= {1'b1, 24'h5851_0a};
      10'd308: {o_verify, o_data} <= {1'b1, 24'h5852_0f};
      10'd309: {o_verify, o_data} <= {1'b1, 24'h5853_0e};
      10'd310: {o_verify, o_data} <= {1'b1, 24'h5854_10};
      10'd311: {o_verify, o_data} <= {1'b1, 24'h5855_10};
      10'd312: {o_verify, o_data} <= {1'b1, 24'h5856_10};
      10'd313: {o_verify, o_data} <= {1'b1, 24'h5857_0a};
      10'd314: {o_verify, o_data} <= {1'b1, 24'h5858_0e};
      10'd315: {o_verify, o_data} <= {1'b1, 24'h5859_0e};
      10'd316: {o_verify, o_data} <= {1'b1, 24'h585a_0f};
      10'd317: {o_verify, o_data} <= {1'b1, 24'h585b_0f};
      10'd318: {o_verify, o_data} <= {1'b1, 24'h585c_0f};
      10'd319: {o_verify, o_data} <= {1'b1, 24'h585d_0a};
      10'd320: {o_verify, o_data} <= {1'b1, 24'h585e_09};
      10'd321: {o_verify, o_data} <= {1'b1, 24'h585f_0d};
      10'd322: {o_verify, o_data} <= {1'b1, 24'h5860_0c};
      10'd323: {o_verify, o_data} <= {1'b1, 24'h5861_0b};
      10'd324: {o_verify, o_data} <= {1'b1, 24'h5862_0d};
      10'd325: {o_verify, o_data} <= {1'b1, 24'h5863_07};
      10'd326: {o_verify, o_data} <= {1'b1, 24'h5864_17};
      10'd327: {o_verify, o_data} <= {1'b1, 24'h5865_14};
      10'd328: {o_verify, o_data} <= {1'b1, 24'h5866_18};
      10'd329: {o_verify, o_data} <= {1'b1, 24'h5867_18};
      10'd330: {o_verify, o_data} <= {1'b1, 24'h5868_16};
      10'd331: {o_verify, o_data} <= {1'b1, 24'h5869_12};
      10'd332: {o_verify, o_data} <= {1'b1, 24'h586a_1b};
      10'd333: {o_verify, o_data} <= {1'b1, 24'h586b_1a};
      10'd334: {o_verify, o_data} <= {1'b1, 24'h586c_16};
      10'd335: {o_verify, o_data} <= {1'b1, 24'h586d_16};
      10'd336: {o_verify, o_data} <= {1'b1, 24'h586e_18};
      10'd337: {o_verify, o_data} <= {1'b1, 24'h586f_1f};
      10'd338: {o_verify, o_data} <= {1'b1, 24'h5870_1c};
      10'd339: {o_verify, o_data} <= {1'b1, 24'h5871_16};
      10'd340: {o_verify, o_data} <= {1'b1, 24'h5872_10};
      10'd341: {o_verify, o_data} <= {1'b1, 24'h5873_0f};
      10'd342: {o_verify, o_data} <= {1'b1, 24'h5874_13};
      10'd343: {o_verify, o_data} <= {1'b1, 24'h5875_1c};
      10'd344: {o_verify, o_data} <= {1'b1, 24'h5876_1e};
      10'd345: {o_verify, o_data} <= {1'b1, 24'h5877_17};
      10'd346: {o_verify, o_data} <= {1'b1, 24'h5878_11};
      10'd347: {o_verify, o_data} <= {1'b1, 24'h5879_11};
      10'd348: {o_verify, o_data} <= {1'b1, 24'h587a_14};
      10'd349: {o_verify, o_data} <= {1'b1, 24'h587b_1e};
      10'd350: {o_verify, o_data} <= {1'b1, 24'h587c_1c};
      10'd351: {o_verify, o_data} <= {1'b1, 24'h587d_1c};
      10'd352: {o_verify, o_data} <= {1'b1, 24'h587e_1a};
      10'd353: {o_verify, o_data} <= {1'b1, 24'h587f_1a};
      10'd354: {o_verify, o_data} <= {1'b1, 24'h5880_1b};
      10'd355: {o_verify, o_data} <= {1'b1, 24'h5881_1f};
      10'd356: {o_verify, o_data} <= {1'b1, 24'h5882_14};
      10'd357: {o_verify, o_data} <= {1'b1, 24'h5883_1a};
      10'd358: {o_verify, o_data} <= {1'b1, 24'h5884_1d};
      10'd359: {o_verify, o_data} <= {1'b1, 24'h5885_1e};
      10'd360: {o_verify, o_data} <= {1'b1, 24'h5886_1a};
      10'd361: {o_verify, o_data} <= {1'b1, 24'h5887_1a};
      10'd362: {o_verify, o_data} <= {1'b1, 24'h5180_ff};
      10'd363: {o_verify, o_data} <= {1'b1, 24'h5181_52};
      10'd364: {o_verify, o_data} <= {1'b1, 24'h5182_11};
      10'd365: {o_verify, o_data} <= {1'b1, 24'h5183_14};
      10'd366: {o_verify, o_data} <= {1'b1, 24'h5184_25};
      10'd367: {o_verify, o_data} <= {1'b1, 24'h5185_24};
      10'd368: {o_verify, o_data} <= {1'b1, 24'h5186_14};
      10'd369: {o_verify, o_data} <= {1'b1, 24'h5187_14};
      10'd370: {o_verify, o_data} <= {1'b1, 24'h5188_14};
      10'd371: {o_verify, o_data} <= {1'b1, 24'h5189_69};
      10'd372: {o_verify, o_data} <= {1'b1, 24'h518a_60};
      10'd373: {o_verify, o_data} <= {1'b1, 24'h518b_a2};
      10'd374: {o_verify, o_data} <= {1'b1, 24'h518c_9c};
      10'd375: {o_verify, o_data} <= {1'b1, 24'h518d_36};
      10'd376: {o_verify, o_data} <= {1'b1, 24'h518e_34};
      10'd377: {o_verify, o_data} <= {1'b1, 24'h518f_54};
      10'd378: {o_verify, o_data} <= {1'b1, 24'h5190_4c};
      10'd379: {o_verify, o_data} <= {1'b1, 24'h5191_f8};
      10'd380: {o_verify, o_data} <= {1'b1, 24'h5192_04};
      10'd381: {o_verify, o_data} <= {1'b1, 24'h5193_70};
      10'd382: {o_verify, o_data} <= {1'b1, 24'h5194_f0};
      10'd383: {o_verify, o_data} <= {1'b1, 24'h5195_f0};
      10'd384: {o_verify, o_data} <= {1'b1, 24'h5196_03};
      10'd385: {o_verify, o_data} <= {1'b1, 24'h5197_01};
      10'd386: {o_verify, o_data} <= {1'b1, 24'h5198_05};
      10'd387: {o_verify, o_data} <= {1'b1, 24'h5199_2f};
      10'd388: {o_verify, o_data} <= {1'b1, 24'h519a_04};
      10'd389: {o_verify, o_data} <= {1'b1, 24'h519b_00};
      10'd390: {o_verify, o_data} <= {1'b1, 24'h519c_06};
      10'd391: {o_verify, o_data} <= {1'b1, 24'h519d_a0};
      10'd392: {o_verify, o_data} <= {1'b1, 24'h519e_a0};
      10'd393: {o_verify, o_data} <= {1'b1, 24'h528a_00};
      10'd394: {o_verify, o_data} <= {1'b1, 24'h528b_01};
      10'd395: {o_verify, o_data} <= {1'b1, 24'h528c_04};
      10'd396: {o_verify, o_data} <= {1'b1, 24'h528d_08};
      10'd397: {o_verify, o_data} <= {1'b1, 24'h528e_10};
      10'd398: {o_verify, o_data} <= {1'b1, 24'h528f_20};
      10'd399: {o_verify, o_data} <= {1'b1, 24'h5290_30};
      10'd400: {o_verify, o_data} <= {1'b1, 24'h5292_00};
      10'd401: {o_verify, o_data} <= {1'b1, 24'h5293_00};
      10'd402: {o_verify, o_data} <= {1'b1, 24'h5294_00};
      10'd403: {o_verify, o_data} <= {1'b1, 24'h5295_01};
      10'd404: {o_verify, o_data} <= {1'b1, 24'h5296_00};
      10'd405: {o_verify, o_data} <= {1'b1, 24'h5297_04};
      10'd406: {o_verify, o_data} <= {1'b1, 24'h5298_00};
      10'd407: {o_verify, o_data} <= {1'b1, 24'h5299_08};
      10'd408: {o_verify, o_data} <= {1'b1, 24'h529a_00};
      10'd409: {o_verify, o_data} <= {1'b1, 24'h529b_10};
      10'd410: {o_verify, o_data} <= {1'b1, 24'h529c_00};
      10'd411: {o_verify, o_data} <= {1'b1, 24'h529d_20};
      10'd412: {o_verify, o_data} <= {1'b1, 24'h529e_00};
      10'd413: {o_verify, o_data} <= {1'b1, 24'h529f_30};
      10'd414: {o_verify, o_data} <= {1'b1, 24'h5282_00};
      10'd415: {o_verify, o_data} <= {1'b1, 24'h5300_00};
      10'd416: {o_verify, o_data} <= {1'b1, 24'h5301_20};
      10'd417: {o_verify, o_data} <= {1'b1, 24'h5302_00};
      10'd418: {o_verify, o_data} <= {1'b1, 24'h5303_7c};
      10'd419: {o_verify, o_data} <= {1'b1, 24'h530c_00};
      10'd420: {o_verify, o_data} <= {1'b1, 24'h530d_10};
      10'd421: {o_verify, o_data} <= {1'b1, 24'h530e_20};
      10'd422: {o_verify, o_data} <= {1'b1, 24'h530f_80};
      10'd423: {o_verify, o_data} <= {1'b1, 24'h5310_20};
      10'd424: {o_verify, o_data} <= {1'b1, 24'h5311_80};
      10'd425: {o_verify, o_data} <= {1'b1, 24'h5308_20};
      10'd426: {o_verify, o_data} <= {1'b1, 24'h5309_40};
      10'd427: {o_verify, o_data} <= {1'b1, 24'h5304_00};
      10'd428: {o_verify, o_data} <= {1'b1, 24'h5305_30};
      10'd429: {o_verify, o_data} <= {1'b1, 24'h5306_00};
      10'd430: {o_verify, o_data} <= {1'b1, 24'h5307_80};
      10'd431: {o_verify, o_data} <= {1'b1, 24'h5314_08};
      10'd432: {o_verify, o_data} <= {1'b1, 24'h5315_20};
      10'd433: {o_verify, o_data} <= {1'b1, 24'h5319_30};
      10'd434: {o_verify, o_data} <= {1'b1, 24'h5316_10};
      10'd435: {o_verify, o_data} <= {1'b1, 24'h5317_00};
      10'd436: {o_verify, o_data} <= {1'b1, 24'h5318_02};
      10'd437: {o_verify, o_data} <= {1'b1, 24'h5380_01};
      10'd438: {o_verify, o_data} <= {1'b1, 24'h5381_00};
      10'd439: {o_verify, o_data} <= {1'b1, 24'h5382_00};
      10'd440: {o_verify, o_data} <= {1'b1, 24'h5383_1f};
      10'd441: {o_verify, o_data} <= {1'b1, 24'h5384_00};
      10'd442: {o_verify, o_data} <= {1'b1, 24'h5385_06};
      10'd443: {o_verify, o_data} <= {1'b1, 24'h5386_00};
      10'd444: {o_verify, o_data} <= {1'b1, 24'h5387_00};
      10'd445: {o_verify, o_data} <= {1'b1, 24'h5388_00};
      10'd446: {o_verify, o_data} <= {1'b1, 24'h5389_e1};
      10'd447: {o_verify, o_data} <= {1'b1, 24'h538a_00};
      10'd448: {o_verify, o_data} <= {1'b1, 24'h538b_2b};
      10'd449: {o_verify, o_data} <= {1'b1, 24'h538c_00};
      10'd450: {o_verify, o_data} <= {1'b1, 24'h538d_00};
      10'd451: {o_verify, o_data} <= {1'b1, 24'h538e_00};
      10'd452: {o_verify, o_data} <= {1'b1, 24'h538f_10};
      10'd453: {o_verify, o_data} <= {1'b1, 24'h5390_00};
      10'd454: {o_verify, o_data} <= {1'b1, 24'h5391_b3};
      10'd455: {o_verify, o_data} <= {1'b1, 24'h5392_00};
      10'd456: {o_verify, o_data} <= {1'b1, 24'h5393_a6};
      10'd457: {o_verify, o_data} <= {1'b1, 24'h5394_08};
      10'd458: {o_verify, o_data} <= {1'b1, 24'h5480_0c};
      10'd459: {o_verify, o_data} <= {1'b1, 24'h5481_18};
      10'd460: {o_verify, o_data} <= {1'b1, 24'h5482_2f};
      10'd461: {o_verify, o_data} <= {1'b1, 24'h5483_55};
      10'd462: {o_verify, o_data} <= {1'b1, 24'h5484_64};
      10'd463: {o_verify, o_data} <= {1'b1, 24'h5485_71};
      10'd464: {o_verify, o_data} <= {1'b1, 24'h5486_7d};
      10'd465: {o_verify, o_data} <= {1'b1, 24'h5487_87};
      10'd466: {o_verify, o_data} <= {1'b1, 24'h5488_91};
      10'd467: {o_verify, o_data} <= {1'b1, 24'h5489_9a};
      10'd468: {o_verify, o_data} <= {1'b1, 24'h548a_aa};
      10'd469: {o_verify, o_data} <= {1'b1, 24'h548b_b8};
      10'd470: {o_verify, o_data} <= {1'b1, 24'h548c_cd};
      10'd471: {o_verify, o_data} <= {1'b1, 24'h548d_dd};
      10'd472: {o_verify, o_data} <= {1'b1, 24'h548e_ea};
      10'd473: {o_verify, o_data} <= {1'b1, 24'h548f_1d};
      10'd474: {o_verify, o_data} <= {1'b1, 24'h5490_05};
      10'd475: {o_verify, o_data} <= {1'b1, 24'h5491_00};
      10'd476: {o_verify, o_data} <= {1'b1, 24'h5492_04};
      10'd477: {o_verify, o_data} <= {1'b1, 24'h5493_20};
      10'd478: {o_verify, o_data} <= {1'b1, 24'h5494_03};
      10'd479: {o_verify, o_data} <= {1'b1, 24'h5495_60};
      10'd480: {o_verify, o_data} <= {1'b1, 24'h5496_02};
      10'd481: {o_verify, o_data} <= {1'b1, 24'h5497_b8};
      10'd482: {o_verify, o_data} <= {1'b1, 24'h5498_02};
      10'd483: {o_verify, o_data} <= {1'b1, 24'h5499_86};
      10'd484: {o_verify, o_data} <= {1'b1, 24'h549a_02};
      10'd485: {o_verify, o_data} <= {1'b1, 24'h549b_5b};
      10'd486: {o_verify, o_data} <= {1'b1, 24'h549c_02};
      10'd487: {o_verify, o_data} <= {1'b1, 24'h549d_3b};
      10'd488: {o_verify, o_data} <= {1'b1, 24'h549e_02};
      10'd489: {o_verify, o_data} <= {1'b1, 24'h549f_1c};
      10'd490: {o_verify, o_data} <= {1'b1, 24'h54a0_02};
      10'd491: {o_verify, o_data} <= {1'b1, 24'h54a1_04};
      10'd492: {o_verify, o_data} <= {1'b1, 24'h54a2_01};
      10'd493: {o_verify, o_data} <= {1'b1, 24'h54a3_ed};
      10'd494: {o_verify, o_data} <= {1'b1, 24'h54a4_01};
      10'd495: {o_verify, o_data} <= {1'b1, 24'h54a5_c5};
      10'd496: {o_verify, o_data} <= {1'b1, 24'h54a6_01};
      10'd497: {o_verify, o_data} <= {1'b1, 24'h54a7_a5};
      10'd498: {o_verify, o_data} <= {1'b1, 24'h54a8_01};
      10'd499: {o_verify, o_data} <= {1'b1, 24'h54a9_6c};
      10'd500: {o_verify, o_data} <= {1'b1, 24'h54aa_01};
      10'd501: {o_verify, o_data} <= {1'b1, 24'h54ab_41};
      10'd502: {o_verify, o_data} <= {1'b1, 24'h54ac_01};
      10'd503: {o_verify, o_data} <= {1'b1, 24'h54ad_20};
      10'd504: {o_verify, o_data} <= {1'b1, 24'h54ae_00};
      10'd505: {o_verify, o_data} <= {1'b1, 24'h54af_16};
      10'd506: {o_verify, o_data} <= {1'b1, 24'h54b0_01};
      10'd507: {o_verify, o_data} <= {1'b1, 24'h54b1_20};
      10'd508: {o_verify, o_data} <= {1'b1, 24'h54b2_00};
      10'd509: {o_verify, o_data} <= {1'b1, 24'h54b3_10};
      10'd510: {o_verify, o_data} <= {1'b1, 24'h54b4_00};
      10'd511: {o_verify, o_data} <= {1'b1, 24'h54b5_f0};
      10'd512: {o_verify, o_data} <= {1'b1, 24'h54b6_00};
      10'd513: {o_verify, o_data} <= {1'b1, 24'h54b7_df};
      10'd514: {o_verify, o_data} <= {1'b1, 24'h5402_3f};
      10'd515: {o_verify, o_data} <= {1'b1, 24'h5403_00};
      10'd516: {o_verify, o_data} <= {1'b1, 24'h5500_10};
      10'd517: {o_verify, o_data} <= {1'b1, 24'h5502_00};
      10'd518: {o_verify, o_data} <= {1'b1, 24'h5503_06};
      10'd519: {o_verify, o_data} <= {1'b1, 24'h5504_00};
      10'd520: {o_verify, o_data} <= {1'b1, 24'h5505_7f};
      10'd521: {o_verify, o_data} <= {1'b1, 24'h5025_80};
      10'd522: {o_verify, o_data} <= {1'b1, 24'h3a0f_30};
      10'd523: {o_verify, o_data} <= {1'b1, 24'h3a10_28};
      10'd524: {o_verify, o_data} <= {1'b1, 24'h3a1b_30};
      10'd525: {o_verify, o_data} <= {1'b1, 24'h3a1e_28};
      10'd526: {o_verify, o_data} <= {1'b1, 24'h3a11_61};
      10'd527: {o_verify, o_data} <= {1'b1, 24'h3a1f_10};
      10'd528: {o_verify, o_data} <= {1'b1, 24'h5688_fd};
      10'd529: {o_verify, o_data} <= {1'b1, 24'h5689_df};
      10'd530: {o_verify, o_data} <= {1'b1, 24'h568a_fe};
      10'd531: {o_verify, o_data} <= {1'b1, 24'h568b_ef};
      10'd532: {o_verify, o_data} <= {1'b1, 24'h568c_fe};
      10'd533: {o_verify, o_data} <= {1'b1, 24'h568d_ef};
      10'd534: {o_verify, o_data} <= {1'b1, 24'h568e_aa};
      10'd535: {o_verify, o_data} <= {1'b1, 24'h568f_aa};*/
      default: {o_verify, o_data} = {1'b0, 24'hffff_ff};
    endcase
  end
    
endmodule